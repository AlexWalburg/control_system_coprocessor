module data_channel
  #(parameter REG_WIDTH 32*12)
   (
    input		  clk,
    input		  rst,
    input		  param_en,
    input [REG_WIDTH-1:0] regs
    );
   
endmodule // data_channel
